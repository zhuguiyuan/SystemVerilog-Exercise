package mlp_pkg;

endpackage